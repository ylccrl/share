`ifndef DMEM_TYPE
`define DMEM_TYPE

`define LD_B    4'b0000
`define LD_H    4'b0001
`define LD_W    4'b0010
`define ST_B    4'b0100
`define ST_H    4'b0101
`define ST_W    4'b0110
`define LD_BU   4'b1000
`define LD_HU   4'b1001

`endif 