`ifndef BR_TYPE
`define BR_TYPE

`define JIRL_B     0011
`define B_B        0100
`define BL_B       0101
`define BEQ_B      0110
`define BNE_B      0111
`define BLT_B      1000
`define BGE_B      1001
`define BLTU_B     1010
`define BGEU_B    1011

`endif