`ifndef BR_TYPE
`define BR_TYPE

`define JIRL_B     4'b0011
`define B_B        4'b0100
`define BL_B       4'b0101
`define BEQ_B      4'b0110
`define BNE_B      4'b0111
`define BLT_B      4'b1000
`define BGE_B      4'b1001
`define BLTU_B     4'b1010
`define BGEU_B     4'b1011

`endif