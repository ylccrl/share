`ifndef BR_TYPE
`define BR_TYPE

`define JIRL_B     6'b010011
`define B_B        6'b010100
`define BL_B       6'b010101
`define BEQ_B      6'b010110
`define BNE_B      6'b010111
`define BLT_B      6'b011000
`define BGE_B      6'b011001
`define BLTU_B     6'b011010
`define BGEU_B     6'b011011

`endif