`ifndef DMEM_TYPE
`define DMEM_TYPE

`define LD_B_D    4'b0000
`define LD_H_D    4'b0001
`define LD_W_D    4'b0010
`define ST_B_D    4'b0100
`define ST_H_D    4'b0101
`define ST_W_D    4'b0110
`define LD_BU_D   4'b1000
`define LD_HU_D   4'b1001

`endif 