module MUX #(
    parameter  WIDTH = 32
    )(
        input   [WIDTH-1:0] src0,src1,
        input   [      0:0] sel,

        output  [WIDTH-1:0] res
    );
    assign res = sel?src1:src0;
endmodule